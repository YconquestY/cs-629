typedef enum {
	Add,
	ShiftL,
	And,
	Not
} InstructionType deriving (Eq,FShow, Bits);

function Bit#(32) alu(InstructionType ins, Bit#(32) v1, Bit#(32) v2);
	return 0;
endfunction

